`timescale 10 ps/10 ps

module DTFM_tb();
reg 				clk = 0;
reg 				clk80 = 0;
reg 				dCLK = 0, dFM = 0, dDAT = 0;
reg	[3:0]		bitCnt	=	15;
reg	[4:0]		wrdCnt	=	19;
reg	[5:0]		strNum	=	63;
reg	[8:0]		frmNum	=	1023;
reg	[9:0]		wrdCnt2	=	1407;

wire				out;


initial begin						// clk ~32768MHz
	clk = 0;
	forever #1525 clk = ~clk;
end

initial begin						// clk ~32768MHz
	clk80 = 0;
	forever #625 clk80 = ~clk80;
end

initial begin						// clk ~1MHz
	dCLK = 0;
	forever #50000 dCLK = ~dCLK;
end

// Static
reg	[11:0]	OK1	=	12'd1101;
reg	[11:0]	OK2	=	12'd1202;
reg	[11:0]	OK3	=	12'd1303;
reg	[11:0]	VK1	=	12'd0;
reg	[11:0]	VK2	=	12'd240;
reg	[11:0]	VK3	=	12'd3855;
reg	[11:0]	UF1	=	12'd1365;
reg	[11:0]	UF2	=	12'd2730;
reg	[11:0]	UF3	=	12'd4095;
reg	[7:0]		corr	=	8'd101;
reg	[7:0]		pel	=	8'd111;
reg	[7:0]		XD		=	8'd121;
reg	[7:0]		YD		=	8'd131;
reg	[7:0]		RM		=	8'd141;
reg	[7:0]		POS	=	8'd151;
reg	[7:0]		ARU	=	8'd161;
// Structure
wire	[15:0]	w[0:1407];
assign w[0] = 16'b0000000000000000; 
assign w[1] = 16'b0000010000000001; 
assign w[2] = 16'b0000000000110000; 
assign w[3] = 16'b0000100000000001; 
assign w[4] = 16'b0100000000110000; 
assign w[5] = 16'b0000011100000001; 
assign w[6] = 16'b0000000000100100; 
assign w[7] = 16'b0000010100000000; 
assign w[8] = 16'b1011000000011000; 
assign w[9] = 16'b0000001101000000; 
assign w[10] = 16'b0111000000001111; 
assign w[11] = 16'b0000001000000000; 
assign w[12] = 16'b0100010000001001; 
assign w[13] = 16'b0000000100110000; 
assign w[14] = 16'b0010100000000101; 
assign w[15] = 16'b0100000010110000; 
assign w[16] = 16'b0001011100000011; 
assign w[17] = 16'b0000000001100100; 
assign w[18] = 16'b0000110100000001; 
assign w[19] = 16'b1011000000111000; 
assign w[20] = 16'b0000011101000000; 
assign w[21] = 16'b1111000000011111; 
assign w[22] = 16'b0000010000000000; 
assign w[23] = 16'b1000010000010001; 
assign w[24] = 16'b0000001000110000; 
assign w[25] = 16'b0100100000001001; 
assign w[26] = 16'b0100000100110000; 
assign w[27] = 16'b0010011100000101; 
assign w[28] = 16'b0000000010100100; 
assign w[29] = 16'b0001010100000010; 
assign w[30] = 16'b1011000001011000; 
assign w[31] = 16'b0000101101000001; 
assign w[32] = 16'b0111000000101111; 
assign w[33] = 16'b0000011000000000; 
assign w[34] = 16'b1100010000011001; 
assign w[35] = 16'b0000001100110000; 
assign w[36] = 16'b0110100000001101; 
assign w[37] = 16'b0100000110110000; 
assign w[38] = 16'b0011011100000111; 
assign w[39] = 16'b0000000011100100; 
assign w[40] = 16'b0001110100000011; 
assign w[41] = 16'b1011000001111000; 
assign w[42] = 16'b0000111101000001; 
assign w[43] = 16'b1111000000111111; 
assign w[44] = 16'b0000100000000001; 
assign w[45] = 16'b0000010000100001; 
assign w[46] = 16'b0000010000110000; 
assign w[47] = 16'b1000100000010001; 
assign w[48] = 16'b0100001000110000; 
assign w[49] = 16'b0100011100001001; 
assign w[50] = 16'b0000000100100100; 
assign w[51] = 16'b0010010100000100; 
assign w[52] = 16'b1011000010011000; 
assign w[53] = 16'b0001001101000010; 
assign w[54] = 16'b0111000001001111; 
assign w[55] = 16'b0000101000000001; 
assign w[56] = 16'b0100010000101001; 
assign w[57] = 16'b0000010100110000; 
assign w[58] = 16'b1010100000010101; 
assign w[59] = 16'b0100001010110000; 
assign w[60] = 16'b0101011100001011; 
assign w[61] = 16'b0000000101100100; 
assign w[62] = 16'b0010110100000101; 
assign w[63] = 16'b1011000010111000; 
assign w[64] = 16'b0001011101000010; 
assign w[65] = 16'b1111000001011111; 
assign w[66] = 16'b0000110000000001; 
assign w[67] = 16'b1000010000110001; 
assign w[68] = 16'b0000011000110000; 
assign w[69] = 16'b1100100000011001; 
assign w[70] = 16'b0100001100110000; 
assign w[71] = 16'b0110011100001101; 
assign w[72] = 16'b0000000110100100; 
assign w[73] = 16'b0011010100000110; 
assign w[74] = 16'b1011000011011000; 
assign w[75] = 16'b0001101101000011; 
assign w[76] = 16'b0111000001101111; 
assign w[77] = 16'b0000111000000001; 
assign w[78] = 16'b1100010000111001; 
assign w[79] = 16'b0000011100110000; 
assign w[80] = 16'b1110100000011101; 
assign w[81] = 16'b0100001110110000; 
assign w[82] = 16'b0111011100001111; 
assign w[83] = 16'b0000000111100100; 
assign w[84] = 16'b0011110100000111; 
assign w[85] = 16'b1011000011111000; 
assign w[86] = 16'b0001111101000011; 
assign w[87] = 16'b1111000001111111; 
assign w[88] = 16'b0001000000000010; 
assign w[89] = 16'b0000010001000001; 
assign w[90] = 16'b0000100000110001; 
assign w[91] = 16'b0000100000100001; 
assign w[92] = 16'b0100010000110000; 
assign w[93] = 16'b1000011100010001; 
assign w[94] = 16'b0000001000100100; 
assign w[95] = 16'b0100010100001000; 
assign w[96] = 16'b1011000100011000; 
assign w[97] = 16'b0010001101000100; 
assign w[98] = 16'b0111000010001111; 
assign w[99] = 16'b0001001000000010; 
assign w[100] = 16'b0100010001001001; 
assign w[101] = 16'b0000100100110001; 
assign w[102] = 16'b0010100000100101; 
assign w[103] = 16'b0100010010110000; 
assign w[104] = 16'b1001011100010011; 
assign w[105] = 16'b0000001001100100; 
assign w[106] = 16'b0100110100001001; 
assign w[107] = 16'b1011000100111000; 
assign w[108] = 16'b0010011101000100; 
assign w[109] = 16'b1111000010011111; 
assign w[110] = 16'b0001010000000010; 
assign w[111] = 16'b1000010001010001; 
assign w[112] = 16'b0000101000110001; 
assign w[113] = 16'b0100100000101001; 
assign w[114] = 16'b0100010100110000; 
assign w[115] = 16'b1010011100010101; 
assign w[116] = 16'b0000001010100100; 
assign w[117] = 16'b0101010100001010; 
assign w[118] = 16'b1011000101011000; 
assign w[119] = 16'b0010101101000101; 
assign w[120] = 16'b0111000010101111; 
assign w[121] = 16'b0001011000000010; 
assign w[122] = 16'b1100010001011001; 
assign w[123] = 16'b0000101100110001; 
assign w[124] = 16'b0110100000101101; 
assign w[125] = 16'b0100010110110000; 
assign w[126] = 16'b1011011100010111; 
assign w[127] = 16'b0000001011100100; 
assign w[128] = 16'b0101110100001011; 
assign w[129] = 16'b1011000101111000; 
assign w[130] = 16'b0010111101000101; 
assign w[131] = 16'b1111000010111111; 
assign w[132] = 16'b0001100000000011; 
assign w[133] = 16'b0000010001100001; 
assign w[134] = 16'b0000110000110001; 
assign w[135] = 16'b1000100000110001; 
assign w[136] = 16'b0100011000110000; 
assign w[137] = 16'b1100011100011001; 
assign w[138] = 16'b0000001100100100; 
assign w[139] = 16'b0110010100001100; 
assign w[140] = 16'b1011000110011000; 
assign w[141] = 16'b0011001101000110; 
assign w[142] = 16'b0111000011001111; 
assign w[143] = 16'b0001101000000011; 
assign w[144] = 16'b0100010001101001; 
assign w[145] = 16'b0000110100110001; 
assign w[146] = 16'b1010100000110101; 
assign w[147] = 16'b0100011010110000; 
assign w[148] = 16'b1101011100011011; 
assign w[149] = 16'b0000001101100100; 
assign w[150] = 16'b0110110100001101; 
assign w[151] = 16'b1011000110111000; 
assign w[152] = 16'b0011011101000110; 
assign w[153] = 16'b1111000011011111; 
assign w[154] = 16'b0001110000000011; 
assign w[155] = 16'b1000010001110001; 
assign w[156] = 16'b0000111000110001; 
assign w[157] = 16'b1100100000111001; 
assign w[158] = 16'b0100011100110000; 
assign w[159] = 16'b1110011100011101; 
assign w[160] = 16'b0000001110100100; 
assign w[161] = 16'b0111010100001110; 
assign w[162] = 16'b1011000111011000; 
assign w[163] = 16'b0011101101000111; 
assign w[164] = 16'b0111000011101111; 
assign w[165] = 16'b0001111000000011; 
assign w[166] = 16'b1100010001111001; 
assign w[167] = 16'b0000111100110001; 
assign w[168] = 16'b1110100000111101; 
assign w[169] = 16'b0100011110110000; 
assign w[170] = 16'b1111011100011111; 
assign w[171] = 16'b0000001111100100; 
assign w[172] = 16'b0111110100001111; 
assign w[173] = 16'b1011000111111000; 
assign w[174] = 16'b0011111101000111; 
assign w[175] = 16'b1111000011111111; 
assign w[176] = 16'b0010000000000100; 
assign w[177] = 16'b0000010010000001; 
assign w[178] = 16'b0001000000110010; 
assign w[179] = 16'b0000100001000001; 
assign w[180] = 16'b0100100000110001; 
assign w[181] = 16'b0000011100100001; 
assign w[182] = 16'b0000010000100100; 
assign w[183] = 16'b1000010100010000; 
assign w[184] = 16'b1011001000011000; 
assign w[185] = 16'b0100001101001000; 
assign w[186] = 16'b0111000100001111; 
assign w[187] = 16'b0010001000000100; 
assign w[188] = 16'b0100010010001001; 
assign w[189] = 16'b0001000100110010; 
assign w[190] = 16'b0010100001000101; 
assign w[191] = 16'b0100100010110001; 
assign w[192] = 16'b0001011100100011; 
assign w[193] = 16'b0000010001100100; 
assign w[194] = 16'b1000110100010001; 
assign w[195] = 16'b1011001000111000; 
assign w[196] = 16'b0100011101001000; 
assign w[197] = 16'b1111000100011111; 
assign w[198] = 16'b0010010000000100; 
assign w[199] = 16'b1000010010010001; 
assign w[200] = 16'b0001001000110010; 
assign w[201] = 16'b0100100001001001; 
assign w[202] = 16'b0100100100110001; 
assign w[203] = 16'b0010011100100101; 
assign w[204] = 16'b0000010010100100; 
assign w[205] = 16'b1001010100010010; 
assign w[206] = 16'b1011001001011000; 
assign w[207] = 16'b0100101101001001; 
assign w[208] = 16'b0111000100101111; 
assign w[209] = 16'b0010011000000100; 
assign w[210] = 16'b1100010010011001; 
assign w[211] = 16'b0001001100110010; 
assign w[212] = 16'b0110100001001101; 
assign w[213] = 16'b0100100110110001; 
assign w[214] = 16'b0011011100100111; 
assign w[215] = 16'b0000010011100100; 
assign w[216] = 16'b1001110100010011; 
assign w[217] = 16'b1011001001111000; 
assign w[218] = 16'b0100111101001001; 
assign w[219] = 16'b1111000100111111; 
assign w[220] = 16'b0010100000000101; 
assign w[221] = 16'b0000010010100001; 
assign w[222] = 16'b0001010000110010; 
assign w[223] = 16'b1000100001010001; 
assign w[224] = 16'b0100101000110001; 
assign w[225] = 16'b0100011100101001; 
assign w[226] = 16'b0000010100100100; 
assign w[227] = 16'b1010010100010100; 
assign w[228] = 16'b1011001010011000; 
assign w[229] = 16'b0101001101001010; 
assign w[230] = 16'b0111000101001111; 
assign w[231] = 16'b0010101000000101; 
assign w[232] = 16'b0100010010101001; 
assign w[233] = 16'b0001010100110010; 
assign w[234] = 16'b1010100001010101; 
assign w[235] = 16'b0100101010110001; 
assign w[236] = 16'b0101011100101011; 
assign w[237] = 16'b0000010101100100; 
assign w[238] = 16'b1010110100010101; 
assign w[239] = 16'b1011001010111000; 
assign w[240] = 16'b0101011101001010; 
assign w[241] = 16'b1111000101011111; 
assign w[242] = 16'b0010110000000101; 
assign w[243] = 16'b1000010010110001; 
assign w[244] = 16'b0001011000110010; 
assign w[245] = 16'b1100100001011001; 
assign w[246] = 16'b0100101100110001; 
assign w[247] = 16'b0110011100101101; 
assign w[248] = 16'b0000010110100100; 
assign w[249] = 16'b1011010100010110; 
assign w[250] = 16'b1011001011011000; 
assign w[251] = 16'b0101101101001011; 
assign w[252] = 16'b0111000101101111; 
assign w[253] = 16'b0010111000000101; 
assign w[254] = 16'b1100010010111001; 
assign w[255] = 16'b0001011100110010; 
assign w[256] = 16'b1110100001011101; 
assign w[257] = 16'b0100101110110001; 
assign w[258] = 16'b0111011100101111; 
assign w[259] = 16'b0000010111100100; 
assign w[260] = 16'b1011110100010111; 
assign w[261] = 16'b1011001011111000; 
assign w[262] = 16'b0101111101001011; 
assign w[263] = 16'b1111000101111111; 
assign w[264] = 16'b0011000000000110; 
assign w[265] = 16'b0000010011000001; 
assign w[266] = 16'b0001100000110011; 
assign w[267] = 16'b0000100001100001; 
assign w[268] = 16'b0100110000110001; 
assign w[269] = 16'b1000011100110001; 
assign w[270] = 16'b0000011000100100; 
assign w[271] = 16'b1100010100011000; 
assign w[272] = 16'b1011001100011000; 
assign w[273] = 16'b0110001101001100; 
assign w[274] = 16'b0111000110001111; 
assign w[275] = 16'b0011001000000110; 
assign w[276] = 16'b0100010011001001; 
assign w[277] = 16'b0001100100110011; 
assign w[278] = 16'b0010100001100101; 
assign w[279] = 16'b0100110010110001; 
assign w[280] = 16'b1001011100110011; 
assign w[281] = 16'b0000011001100100; 
assign w[282] = 16'b1100110100011001; 
assign w[283] = 16'b1011001100111000; 
assign w[284] = 16'b0110011101001100; 
assign w[285] = 16'b1111000110011111; 
assign w[286] = 16'b0011010000000110; 
assign w[287] = 16'b1000010011010001; 
assign w[288] = 16'b0001101000110011; 
assign w[289] = 16'b0100100001101001; 
assign w[290] = 16'b0100110100110001; 
assign w[291] = 16'b1010011100110101; 
assign w[292] = 16'b0000011010100100; 
assign w[293] = 16'b1101010100011010; 
assign w[294] = 16'b1011001101011000; 
assign w[295] = 16'b0110101101001101; 
assign w[296] = 16'b0111000110101111; 
assign w[297] = 16'b0011011000000110; 
assign w[298] = 16'b1100010011011001; 
assign w[299] = 16'b0001101100110011; 
assign w[300] = 16'b0110100001101101; 
assign w[301] = 16'b0100110110110001; 
assign w[302] = 16'b1011011100110111; 
assign w[303] = 16'b0000011011100100; 
assign w[304] = 16'b1101110100011011; 
assign w[305] = 16'b1011001101111000; 
assign w[306] = 16'b0110111101001101; 
assign w[307] = 16'b1111000110111111; 
assign w[308] = 16'b0011100000000111; 
assign w[309] = 16'b0000010011100001; 
assign w[310] = 16'b0001110000110011; 
assign w[311] = 16'b1000100001110001; 
assign w[312] = 16'b0100111000110001; 
assign w[313] = 16'b1100011100111001; 
assign w[314] = 16'b0000011100100100; 
assign w[315] = 16'b1110010100011100; 
assign w[316] = 16'b1011001110011000; 
assign w[317] = 16'b0111001101001110; 
assign w[318] = 16'b0111000111001111; 
assign w[319] = 16'b0011101000000111; 
assign w[320] = 16'b0100010011101001; 
assign w[321] = 16'b0001110100110011; 
assign w[322] = 16'b1010100001110101; 
assign w[323] = 16'b0100111010110001; 
assign w[324] = 16'b1101011100111011; 
assign w[325] = 16'b0000011101100100; 
assign w[326] = 16'b1110110100011101; 
assign w[327] = 16'b1011001110111000; 
assign w[328] = 16'b0111011101001110; 
assign w[329] = 16'b1111000111011111; 
assign w[330] = 16'b0011110000000111; 
assign w[331] = 16'b1000010011110001; 
assign w[332] = 16'b0001111000110011; 
assign w[333] = 16'b1100100001111001; 
assign w[334] = 16'b0100111100110001; 
assign w[335] = 16'b1110011100111101; 
assign w[336] = 16'b0000011110100100; 
assign w[337] = 16'b1111010100011110; 
assign w[338] = 16'b1011001111011000; 
assign w[339] = 16'b0111101101001111; 
assign w[340] = 16'b0111000111101111; 
assign w[341] = 16'b0011111000000111; 
assign w[342] = 16'b1100010011111001; 
assign w[343] = 16'b0001111100110011; 
assign w[344] = 16'b1110100001111101; 
assign w[345] = 16'b0100111110110001; 
assign w[346] = 16'b1111011100111111; 
assign w[347] = 16'b0000011111100100; 
assign w[348] = 16'b1111110100011111; 
assign w[349] = 16'b1011001111111000; 
assign w[350] = 16'b0111111101001111; 
assign w[351] = 16'b1111000111111111; 
assign w[352] = 16'b0100000000001000; 
assign w[353] = 16'b0000010100000001; 
assign w[354] = 16'b0010000000110100; 
assign w[355] = 16'b0000100010000001; 
assign w[356] = 16'b0101000000110010; 
assign w[357] = 16'b0000011101000001; 
assign w[358] = 16'b0000100000100101; 
assign w[359] = 16'b0000010100100000; 
assign w[360] = 16'b1011010000011000; 
assign w[361] = 16'b1000001101010000; 
assign w[362] = 16'b0111001000001111; 
assign w[363] = 16'b0100001000001000; 
assign w[364] = 16'b0100010100001001; 
assign w[365] = 16'b0010000100110100; 
assign w[366] = 16'b0010100010000101; 
assign w[367] = 16'b0101000010110010; 
assign w[368] = 16'b0001011101000011; 
assign w[369] = 16'b0000100001100101; 
assign w[370] = 16'b0000110100100001; 
assign w[371] = 16'b1011010000111000; 
assign w[372] = 16'b1000011101010000; 
assign w[373] = 16'b1111001000011111; 
assign w[374] = 16'b0100010000001000; 
assign w[375] = 16'b1000010100010001; 
assign w[376] = 16'b0010001000110100; 
assign w[377] = 16'b0100100010001001; 
assign w[378] = 16'b0101000100110010; 
assign w[379] = 16'b0010011101000101; 
assign w[380] = 16'b0000100010100101; 
assign w[381] = 16'b0001010100100010; 
assign w[382] = 16'b1011010001011000; 
assign w[383] = 16'b1000101101010001; 
assign w[384] = 16'b0111001000101111; 
assign w[385] = 16'b0100011000001000; 
assign w[386] = 16'b1100010100011001; 
assign w[387] = 16'b0010001100110100; 
assign w[388] = 16'b0110100010001101; 
assign w[389] = 16'b0101000110110010; 
assign w[390] = 16'b0011011101000111; 
assign w[391] = 16'b0000100011100101; 
assign w[392] = 16'b0001110100100011; 
assign w[393] = 16'b1011010001111000; 
assign w[394] = 16'b1000111101010001; 
assign w[395] = 16'b1111001000111111; 
assign w[396] = 16'b0100100000001001; 
assign w[397] = 16'b0000010100100001; 
assign w[398] = 16'b0010010000110100; 
assign w[399] = 16'b1000100010010001; 
assign w[400] = 16'b0101001000110010; 
assign w[401] = 16'b0100011101001001; 
assign w[402] = 16'b0000100100100101; 
assign w[403] = 16'b0010010100100100; 
assign w[404] = 16'b1011010010011000; 
assign w[405] = 16'b1001001101010010; 
assign w[406] = 16'b0111001001001111; 
assign w[407] = 16'b0100101000001001; 
assign w[408] = 16'b0100010100101001; 
assign w[409] = 16'b0010010100110100; 
assign w[410] = 16'b1010100010010101; 
assign w[411] = 16'b0101001010110010; 
assign w[412] = 16'b0101011101001011; 
assign w[413] = 16'b0000100101100101; 
assign w[414] = 16'b0010110100100101; 
assign w[415] = 16'b1011010010111000; 
assign w[416] = 16'b1001011101010010; 
assign w[417] = 16'b1111001001011111; 
assign w[418] = 16'b0100110000001001; 
assign w[419] = 16'b1000010100110001; 
assign w[420] = 16'b0010011000110100; 
assign w[421] = 16'b1100100010011001; 
assign w[422] = 16'b0101001100110010; 
assign w[423] = 16'b0110011101001101; 
assign w[424] = 16'b0000100110100101; 
assign w[425] = 16'b0011010100100110; 
assign w[426] = 16'b1011010011011000; 
assign w[427] = 16'b1001101101010011; 
assign w[428] = 16'b0111001001101111; 
assign w[429] = 16'b0100111000001001; 
assign w[430] = 16'b1100010100111001; 
assign w[431] = 16'b0010011100110100; 
assign w[432] = 16'b1110100010011101; 
assign w[433] = 16'b0101001110110010; 
assign w[434] = 16'b0111011101001111; 
assign w[435] = 16'b0000100111100101; 
assign w[436] = 16'b0011110100100111; 
assign w[437] = 16'b1011010011111000; 
assign w[438] = 16'b1001111101010011; 
assign w[439] = 16'b1111001001111111; 
assign w[440] = 16'b0101000000001010; 
assign w[441] = 16'b0000010101000001; 
assign w[442] = 16'b0010100000110101; 
assign w[443] = 16'b0000100010100001; 
assign w[444] = 16'b0101010000110010; 
assign w[445] = 16'b1000011101010001; 
assign w[446] = 16'b0000101000100101; 
assign w[447] = 16'b0100010100101000; 
assign w[448] = 16'b1011010100011000; 
assign w[449] = 16'b1010001101010100; 
assign w[450] = 16'b0111001010001111; 
assign w[451] = 16'b0101001000001010; 
assign w[452] = 16'b0100010101001001; 
assign w[453] = 16'b0010100100110101; 
assign w[454] = 16'b0010100010100101; 
assign w[455] = 16'b0101010010110010; 
assign w[456] = 16'b1001011101010011; 
assign w[457] = 16'b0000101001100101; 
assign w[458] = 16'b0100110100101001; 
assign w[459] = 16'b1011010100111000; 
assign w[460] = 16'b1010011101010100; 
assign w[461] = 16'b1111001010011111; 
assign w[462] = 16'b0101010000001010; 
assign w[463] = 16'b1000010101010001; 
assign w[464] = 16'b0010101000110101; 
assign w[465] = 16'b0100100010101001; 
assign w[466] = 16'b0101010100110010; 
assign w[467] = 16'b1010011101010101; 
assign w[468] = 16'b0000101010100101; 
assign w[469] = 16'b0101010100101010; 
assign w[470] = 16'b1011010101011000; 
assign w[471] = 16'b1010101101010101; 
assign w[472] = 16'b0111001010101111; 
assign w[473] = 16'b0101011000001010; 
assign w[474] = 16'b1100010101011001; 
assign w[475] = 16'b0010101100110101; 
assign w[476] = 16'b0110100010101101; 
assign w[477] = 16'b0101010110110010; 
assign w[478] = 16'b1011011101010111; 
assign w[479] = 16'b0000101011100101; 
assign w[480] = 16'b0101110100101011; 
assign w[481] = 16'b1011010101111000; 
assign w[482] = 16'b1010111101010101; 
assign w[483] = 16'b1111001010111111; 
assign w[484] = 16'b0101100000001011; 
assign w[485] = 16'b0000010101100001; 
assign w[486] = 16'b0010110000110101; 
assign w[487] = 16'b1000100010110001; 
assign w[488] = 16'b0101011000110010; 
assign w[489] = 16'b1100011101011001; 
assign w[490] = 16'b0000101100100101; 
assign w[491] = 16'b0110010100101100; 
assign w[492] = 16'b1011010110011000; 
assign w[493] = 16'b1011001101010110; 
assign w[494] = 16'b0111001011001111; 
assign w[495] = 16'b0101101000001011; 
assign w[496] = 16'b0100010101101001; 
assign w[497] = 16'b0010110100110101; 
assign w[498] = 16'b1010100010110101; 
assign w[499] = 16'b0101011010110010; 
assign w[500] = 16'b1101011101011011; 
assign w[501] = 16'b0000101101100101; 
assign w[502] = 16'b0110110100101101; 
assign w[503] = 16'b1011010110111000; 
assign w[504] = 16'b1011011101010110; 
assign w[505] = 16'b1111001011011111; 
assign w[506] = 16'b0101110000001011; 
assign w[507] = 16'b1000010101110001; 
assign w[508] = 16'b0010111000110101; 
assign w[509] = 16'b1100100010111001; 
assign w[510] = 16'b0101011100110010; 
assign w[511] = 16'b1110011101011101; 
assign w[512] = 16'b0000101110100101; 
assign w[513] = 16'b0111010100101110; 
assign w[514] = 16'b1011010111011000; 
assign w[515] = 16'b1011101101010111; 
assign w[516] = 16'b0111001011101111; 
assign w[517] = 16'b0101111000001011; 
assign w[518] = 16'b1100010101111001; 
assign w[519] = 16'b0010111100110101; 
assign w[520] = 16'b1110100010111101; 
assign w[521] = 16'b0101011110110010; 
assign w[522] = 16'b1111011101011111; 
assign w[523] = 16'b0000101111100101; 
assign w[524] = 16'b0111110100101111; 
assign w[525] = 16'b1011010111111000; 
assign w[526] = 16'b1011111101010111; 
assign w[527] = 16'b1111001011111111; 
assign w[528] = 16'b0110000000001100; 
assign w[529] = 16'b0000010110000001; 
assign w[530] = 16'b0011000000110110; 
assign w[531] = 16'b0000100011000001; 
assign w[532] = 16'b0101100000110011; 
assign w[533] = 16'b0000011101100001; 
assign w[534] = 16'b0000110000100101; 
assign w[535] = 16'b1000010100110000; 
assign w[536] = 16'b1011011000011000; 
assign w[537] = 16'b1100001101011000; 
assign w[538] = 16'b0111001100001111; 
assign w[539] = 16'b0110001000001100; 
assign w[540] = 16'b0100010110001001; 
assign w[541] = 16'b0011000100110110; 
assign w[542] = 16'b0010100011000101; 
assign w[543] = 16'b0101100010110011; 
assign w[544] = 16'b0001011101100011; 
assign w[545] = 16'b0000110001100101; 
assign w[546] = 16'b1000110100110001; 
assign w[547] = 16'b1011011000111000; 
assign w[548] = 16'b1100011101011000; 
assign w[549] = 16'b1111001100011111; 
assign w[550] = 16'b0110010000001100; 
assign w[551] = 16'b1000010110010001; 
assign w[552] = 16'b0011001000110110; 
assign w[553] = 16'b0100100011001001; 
assign w[554] = 16'b0101100100110011; 
assign w[555] = 16'b0010011101100101; 
assign w[556] = 16'b0000110010100101; 
assign w[557] = 16'b1001010100110010; 
assign w[558] = 16'b1011011001011000; 
assign w[559] = 16'b1100101101011001; 
assign w[560] = 16'b0111001100101111; 
assign w[561] = 16'b0110011000001100; 
assign w[562] = 16'b1100010110011001; 
assign w[563] = 16'b0011001100110110; 
assign w[564] = 16'b0110100011001101; 
assign w[565] = 16'b0101100110110011; 
assign w[566] = 16'b0011011101100111; 
assign w[567] = 16'b0000110011100101; 
assign w[568] = 16'b1001110100110011; 
assign w[569] = 16'b1011011001111000; 
assign w[570] = 16'b1100111101011001; 
assign w[571] = 16'b1111001100111111; 
assign w[572] = 16'b0110100000001101; 
assign w[573] = 16'b0000010110100001; 
assign w[574] = 16'b0011010000110110; 
assign w[575] = 16'b1000100011010001; 
assign w[576] = 16'b0101101000110011; 
assign w[577] = 16'b0100011101101001; 
assign w[578] = 16'b0000110100100101; 
assign w[579] = 16'b1010010100110100; 
assign w[580] = 16'b1011011010011000; 
assign w[581] = 16'b1101001101011010; 
assign w[582] = 16'b0111001101001111; 
assign w[583] = 16'b0110101000001101; 
assign w[584] = 16'b0100010110101001; 
assign w[585] = 16'b0011010100110110; 
assign w[586] = 16'b1010100011010101; 
assign w[587] = 16'b0101101010110011; 
assign w[588] = 16'b0101011101101011; 
assign w[589] = 16'b0000110101100101; 
assign w[590] = 16'b1010110100110101; 
assign w[591] = 16'b1011011010111000; 
assign w[592] = 16'b1101011101011010; 
assign w[593] = 16'b1111001101011111; 
assign w[594] = 16'b0110110000001101; 
assign w[595] = 16'b1000010110110001; 
assign w[596] = 16'b0011011000110110; 
assign w[597] = 16'b1100100011011001; 
assign w[598] = 16'b0101101100110011; 
assign w[599] = 16'b0110011101101101; 
assign w[600] = 16'b0000110110100101; 
assign w[601] = 16'b1011010100110110; 
assign w[602] = 16'b1011011011011000; 
assign w[603] = 16'b1101101101011011; 
assign w[604] = 16'b0111001101101111; 
assign w[605] = 16'b0110111000001101; 
assign w[606] = 16'b1100010110111001; 
assign w[607] = 16'b0011011100110110; 
assign w[608] = 16'b1110100011011101; 
assign w[609] = 16'b0101101110110011; 
assign w[610] = 16'b0111011101101111; 
assign w[611] = 16'b0000110111100101; 
assign w[612] = 16'b1011110100110111; 
assign w[613] = 16'b1011011011111000; 
assign w[614] = 16'b1101111101011011; 
assign w[615] = 16'b1111001101111111; 
assign w[616] = 16'b0111000000001110; 
assign w[617] = 16'b0000010111000001; 
assign w[618] = 16'b0011100000110111; 
assign w[619] = 16'b0000100011100001; 
assign w[620] = 16'b0101110000110011; 
assign w[621] = 16'b1000011101110001; 
assign w[622] = 16'b0000111000100101; 
assign w[623] = 16'b1100010100111000; 
assign w[624] = 16'b1011011100011000; 
assign w[625] = 16'b1110001101011100; 
assign w[626] = 16'b0111001110001111; 
assign w[627] = 16'b0111001000001110; 
assign w[628] = 16'b0100010111001001; 
assign w[629] = 16'b0011100100110111; 
assign w[630] = 16'b0010100011100101; 
assign w[631] = 16'b0101110010110011; 
assign w[632] = 16'b1001011101110011; 
assign w[633] = 16'b0000111001100101; 
assign w[634] = 16'b1100110100111001; 
assign w[635] = 16'b1011011100111000; 
assign w[636] = 16'b1110011101011100; 
assign w[637] = 16'b1111001110011111; 
assign w[638] = 16'b0111010000001110; 
assign w[639] = 16'b1000010111010001; 
assign w[640] = 16'b0011101000110111; 
assign w[641] = 16'b0100100011101001; 
assign w[642] = 16'b0101110100110011; 
assign w[643] = 16'b1010011101110101; 
assign w[644] = 16'b0000111010100101; 
assign w[645] = 16'b1101010100111010; 
assign w[646] = 16'b1011011101011000; 
assign w[647] = 16'b1110101101011101; 
assign w[648] = 16'b0111001110101111; 
assign w[649] = 16'b0111011000001110; 
assign w[650] = 16'b1100010111011001; 
assign w[651] = 16'b0011101100110111; 
assign w[652] = 16'b0110100011101101; 
assign w[653] = 16'b0101110110110011; 
assign w[654] = 16'b1011011101110111; 
assign w[655] = 16'b0000111011100101; 
assign w[656] = 16'b1101110100111011; 
assign w[657] = 16'b1011011101111000; 
assign w[658] = 16'b1110111101011101; 
assign w[659] = 16'b1111001110111111; 
assign w[660] = 16'b0111100000001111; 
assign w[661] = 16'b0000010111100001; 
assign w[662] = 16'b0011110000110111; 
assign w[663] = 16'b1000100011110001; 
assign w[664] = 16'b0101111000110011; 
assign w[665] = 16'b1100011101111001; 
assign w[666] = 16'b0000111100100101; 
assign w[667] = 16'b1110010100111100; 
assign w[668] = 16'b1011011110011000; 
assign w[669] = 16'b1111001101011110; 
assign w[670] = 16'b0111001111001111; 
assign w[671] = 16'b0111101000001111; 
assign w[672] = 16'b0100010111101001; 
assign w[673] = 16'b0011110100110111; 
assign w[674] = 16'b1010100011110101; 
assign w[675] = 16'b0101111010110011; 
assign w[676] = 16'b1101011101111011; 
assign w[677] = 16'b0000111101100101; 
assign w[678] = 16'b1110110100111101; 
assign w[679] = 16'b1011011110111000; 
assign w[680] = 16'b1111011101011110; 
assign w[681] = 16'b1111001111011111; 
assign w[682] = 16'b0111110000001111; 
assign w[683] = 16'b1000010111110001; 
assign w[684] = 16'b0011111000110111; 
assign w[685] = 16'b1100100011111001; 
assign w[686] = 16'b0101111100110011; 
assign w[687] = 16'b1110011101111101; 
assign w[688] = 16'b0000111110100101; 
assign w[689] = 16'b1111010100111110; 
assign w[690] = 16'b1011011111011000; 
assign w[691] = 16'b1111101101011111; 
assign w[692] = 16'b0111001111101111; 
assign w[693] = 16'b0111111000001111; 
assign w[694] = 16'b1100010111111001; 
assign w[695] = 16'b0011111100110111; 
assign w[696] = 16'b1110100011111101; 
assign w[697] = 16'b0101111110110011; 
assign w[698] = 16'b1111011101111111; 
assign w[699] = 16'b0000111111100101; 
assign w[700] = 16'b1111110100111111; 
assign w[701] = 16'b1011011111111000; 
assign w[702] = 16'b1111111101011111; 
assign w[703] = 16'b1111001111111111; 
assign w[704] = 16'b1000000000010000; 
assign w[705] = 16'b0000011000000001; 
assign w[706] = 16'b0100000000111000; 
assign w[707] = 16'b0000100100000001; 
assign w[708] = 16'b0110000000110100; 
assign w[709] = 16'b0000011110000001; 
assign w[710] = 16'b0001000000100110; 
assign w[711] = 16'b0000010101000000; 
assign w[712] = 16'b1011100000011001; 
assign w[713] = 16'b0000001101100000; 
assign w[714] = 16'b0111010000001111; 
assign w[715] = 16'b1000001000010000; 
assign w[716] = 16'b0100011000001001; 
assign w[717] = 16'b0100000100111000; 
assign w[718] = 16'b0010100100000101; 
assign w[719] = 16'b0110000010110100; 
assign w[720] = 16'b0001011110000011; 
assign w[721] = 16'b0001000001100110; 
assign w[722] = 16'b0000110101000001; 
assign w[723] = 16'b1011100000111001; 
assign w[724] = 16'b0000011101100000; 
assign w[725] = 16'b1111010000011111; 
assign w[726] = 16'b1000010000010000; 
assign w[727] = 16'b1000011000010001; 
assign w[728] = 16'b0100001000111000; 
assign w[729] = 16'b0100100100001001; 
assign w[730] = 16'b0110000100110100; 
assign w[731] = 16'b0010011110000101; 
assign w[732] = 16'b0001000010100110; 
assign w[733] = 16'b0001010101000010; 
assign w[734] = 16'b1011100001011001; 
assign w[735] = 16'b0000101101100001; 
assign w[736] = 16'b0111010000101111; 
assign w[737] = 16'b1000011000010000; 
assign w[738] = 16'b1100011000011001; 
assign w[739] = 16'b0100001100111000; 
assign w[740] = 16'b0110100100001101; 
assign w[741] = 16'b0110000110110100; 
assign w[742] = 16'b0011011110000111; 
assign w[743] = 16'b0001000011100110; 
assign w[744] = 16'b0001110101000011; 
assign w[745] = 16'b1011100001111001; 
assign w[746] = 16'b0000111101100001; 
assign w[747] = 16'b1111010000111111; 
assign w[748] = 16'b1000100000010001; 
assign w[749] = 16'b0000011000100001; 
assign w[750] = 16'b0100010000111000; 
assign w[751] = 16'b1000100100010001; 
assign w[752] = 16'b0110001000110100; 
assign w[753] = 16'b0100011110001001; 
assign w[754] = 16'b0001000100100110; 
assign w[755] = 16'b0010010101000100; 
assign w[756] = 16'b1011100010011001; 
assign w[757] = 16'b0001001101100010; 
assign w[758] = 16'b0111010001001111; 
assign w[759] = 16'b1000101000010001; 
assign w[760] = 16'b0100011000101001; 
assign w[761] = 16'b0100010100111000; 
assign w[762] = 16'b1010100100010101; 
assign w[763] = 16'b0110001010110100; 
assign w[764] = 16'b0101011110001011; 
assign w[765] = 16'b0001000101100110; 
assign w[766] = 16'b0010110101000101; 
assign w[767] = 16'b1011100010111001; 
assign w[768] = 16'b0001011101100010; 
assign w[769] = 16'b1111010001011111; 
assign w[770] = 16'b1000110000010001; 
assign w[771] = 16'b1000011000110001; 
assign w[772] = 16'b0100011000111000; 
assign w[773] = 16'b1100100100011001; 
assign w[774] = 16'b0110001100110100; 
assign w[775] = 16'b0110011110001101; 
assign w[776] = 16'b0001000110100110; 
assign w[777] = 16'b0011010101000110; 
assign w[778] = 16'b1011100011011001; 
assign w[779] = 16'b0001101101100011; 
assign w[780] = 16'b0111010001101111; 
assign w[781] = 16'b1000111000010001; 
assign w[782] = 16'b1100011000111001; 
assign w[783] = 16'b0100011100111000; 
assign w[784] = 16'b1110100100011101; 
assign w[785] = 16'b0110001110110100; 
assign w[786] = 16'b0111011110001111; 
assign w[787] = 16'b0001000111100110; 
assign w[788] = 16'b0011110101000111; 
assign w[789] = 16'b1011100011111001; 
assign w[790] = 16'b0001111101100011; 
assign w[791] = 16'b1111010001111111; 
assign w[792] = 16'b1001000000010010; 
assign w[793] = 16'b0000011001000001; 
assign w[794] = 16'b0100100000111001; 
assign w[795] = 16'b0000100100100001; 
assign w[796] = 16'b0110010000110100; 
assign w[797] = 16'b1000011110010001; 
assign w[798] = 16'b0001001000100110; 
assign w[799] = 16'b0100010101001000; 
assign w[800] = 16'b1011100100011001; 
assign w[801] = 16'b0010001101100100; 
assign w[802] = 16'b0111010010001111; 
assign w[803] = 16'b1001001000010010; 
assign w[804] = 16'b0100011001001001; 
assign w[805] = 16'b0100100100111001; 
assign w[806] = 16'b0010100100100101; 
assign w[807] = 16'b0110010010110100; 
assign w[808] = 16'b1001011110010011; 
assign w[809] = 16'b0001001001100110; 
assign w[810] = 16'b0100110101001001; 
assign w[811] = 16'b1011100100111001; 
assign w[812] = 16'b0010011101100100; 
assign w[813] = 16'b1111010010011111; 
assign w[814] = 16'b1001010000010010; 
assign w[815] = 16'b1000011001010001; 
assign w[816] = 16'b0100101000111001; 
assign w[817] = 16'b0100100100101001; 
assign w[818] = 16'b0110010100110100; 
assign w[819] = 16'b1010011110010101; 
assign w[820] = 16'b0001001010100110; 
assign w[821] = 16'b0101010101001010; 
assign w[822] = 16'b1011100101011001; 
assign w[823] = 16'b0010101101100101; 
assign w[824] = 16'b0111010010101111; 
assign w[825] = 16'b1001011000010010; 
assign w[826] = 16'b1100011001011001; 
assign w[827] = 16'b0100101100111001; 
assign w[828] = 16'b0110100100101101; 
assign w[829] = 16'b0110010110110100; 
assign w[830] = 16'b1011011110010111; 
assign w[831] = 16'b0001001011100110; 
assign w[832] = 16'b0101110101001011; 
assign w[833] = 16'b1011100101111001; 
assign w[834] = 16'b0010111101100101; 
assign w[835] = 16'b1111010010111111; 
assign w[836] = 16'b1001100000010011; 
assign w[837] = 16'b0000011001100001; 
assign w[838] = 16'b0100110000111001; 
assign w[839] = 16'b1000100100110001; 
assign w[840] = 16'b0110011000110100; 
assign w[841] = 16'b1100011110011001; 
assign w[842] = 16'b0001001100100110; 
assign w[843] = 16'b0110010101001100; 
assign w[844] = 16'b1011100110011001; 
assign w[845] = 16'b0011001101100110; 
assign w[846] = 16'b0111010011001111; 
assign w[847] = 16'b1001101000010011; 
assign w[848] = 16'b0100011001101001; 
assign w[849] = 16'b0100110100111001; 
assign w[850] = 16'b1010100100110101; 
assign w[851] = 16'b0110011010110100; 
assign w[852] = 16'b1101011110011011; 
assign w[853] = 16'b0001001101100110; 
assign w[854] = 16'b0110110101001101; 
assign w[855] = 16'b1011100110111001; 
assign w[856] = 16'b0011011101100110; 
assign w[857] = 16'b1111010011011111; 
assign w[858] = 16'b1001110000010011; 
assign w[859] = 16'b1000011001110001; 
assign w[860] = 16'b0100111000111001; 
assign w[861] = 16'b1100100100111001; 
assign w[862] = 16'b0110011100110100; 
assign w[863] = 16'b1110011110011101; 
assign w[864] = 16'b0001001110100110; 
assign w[865] = 16'b0111010101001110; 
assign w[866] = 16'b1011100111011001; 
assign w[867] = 16'b0011101101100111; 
assign w[868] = 16'b0111010011101111; 
assign w[869] = 16'b1001111000010011; 
assign w[870] = 16'b1100011001111001; 
assign w[871] = 16'b0100111100111001; 
assign w[872] = 16'b1110100100111101; 
assign w[873] = 16'b0110011110110100; 
assign w[874] = 16'b1111011110011111; 
assign w[875] = 16'b0001001111100110; 
assign w[876] = 16'b0111110101001111; 
assign w[877] = 16'b1011100111111001; 
assign w[878] = 16'b0011111101100111; 
assign w[879] = 16'b1111010011111111; 
assign w[880] = 16'b1010000000010100; 
assign w[881] = 16'b0000011010000001; 
assign w[882] = 16'b0101000000111010; 
assign w[883] = 16'b0000100101000001; 
assign w[884] = 16'b0110100000110101; 
assign w[885] = 16'b0000011110100001; 
assign w[886] = 16'b0001010000100110; 
assign w[887] = 16'b1000010101010000; 
assign w[888] = 16'b1011101000011001; 
assign w[889] = 16'b0100001101101000; 
assign w[890] = 16'b0111010100001111; 
assign w[891] = 16'b1010001000010100; 
assign w[892] = 16'b0100011010001001; 
assign w[893] = 16'b0101000100111010; 
assign w[894] = 16'b0010100101000101; 
assign w[895] = 16'b0110100010110101; 
assign w[896] = 16'b0001011110100011; 
assign w[897] = 16'b0001010001100110; 
assign w[898] = 16'b1000110101010001; 
assign w[899] = 16'b1011101000111001; 
assign w[900] = 16'b0100011101101000; 
assign w[901] = 16'b1111010100011111; 
assign w[902] = 16'b1010010000010100; 
assign w[903] = 16'b1000011010010001; 
assign w[904] = 16'b0101001000111010; 
assign w[905] = 16'b0100100101001001; 
assign w[906] = 16'b0110100100110101; 
assign w[907] = 16'b0010011110100101; 
assign w[908] = 16'b0001010010100110; 
assign w[909] = 16'b1001010101010010; 
assign w[910] = 16'b1011101001011001; 
assign w[911] = 16'b0100101101101001; 
assign w[912] = 16'b0111010100101111; 
assign w[913] = 16'b1010011000010100; 
assign w[914] = 16'b1100011010011001; 
assign w[915] = 16'b0101001100111010; 
assign w[916] = 16'b0110100101001101; 
assign w[917] = 16'b0110100110110101; 
assign w[918] = 16'b0011011110100111; 
assign w[919] = 16'b0001010011100110; 
assign w[920] = 16'b1001110101010011; 
assign w[921] = 16'b1011101001111001; 
assign w[922] = 16'b0100111101101001; 
assign w[923] = 16'b1111010100111111; 
assign w[924] = 16'b1010100000010101; 
assign w[925] = 16'b0000011010100001; 
assign w[926] = 16'b0101010000111010; 
assign w[927] = 16'b1000100101010001; 
assign w[928] = 16'b0110101000110101; 
assign w[929] = 16'b0100011110101001; 
assign w[930] = 16'b0001010100100110; 
assign w[931] = 16'b1010010101010100; 
assign w[932] = 16'b1011101010011001; 
assign w[933] = 16'b0101001101101010; 
assign w[934] = 16'b0111010101001111; 
assign w[935] = 16'b1010101000010101; 
assign w[936] = 16'b0100011010101001; 
assign w[937] = 16'b0101010100111010; 
assign w[938] = 16'b1010100101010101; 
assign w[939] = 16'b0110101010110101; 
assign w[940] = 16'b0101011110101011; 
assign w[941] = 16'b0001010101100110; 
assign w[942] = 16'b1010110101010101; 
assign w[943] = 16'b1011101010111001; 
assign w[944] = 16'b0101011101101010; 
assign w[945] = 16'b1111010101011111; 
assign w[946] = 16'b1010110000010101; 
assign w[947] = 16'b1000011010110001; 
assign w[948] = 16'b0101011000111010; 
assign w[949] = 16'b1100100101011001; 
assign w[950] = 16'b0110101100110101; 
assign w[951] = 16'b0110011110101101; 
assign w[952] = 16'b0001010110100110; 
assign w[953] = 16'b1011010101010110; 
assign w[954] = 16'b1011101011011001; 
assign w[955] = 16'b0101101101101011; 
assign w[956] = 16'b0111010101101111; 
assign w[957] = 16'b1010111000010101; 
assign w[958] = 16'b1100011010111001; 
assign w[959] = 16'b0101011100111010; 
assign w[960] = 16'b1110100101011101; 
assign w[961] = 16'b0110101110110101; 
assign w[962] = 16'b0111011110101111; 
assign w[963] = 16'b0001010111100110; 
assign w[964] = 16'b1011110101010111; 
assign w[965] = 16'b1011101011111001; 
assign w[966] = 16'b0101111101101011; 
assign w[967] = 16'b1111010101111111; 
assign w[968] = 16'b1011000000010110; 
assign w[969] = 16'b0000011011000001; 
assign w[970] = 16'b0101100000111011; 
assign w[971] = 16'b0000100101100001; 
assign w[972] = 16'b0110110000110101; 
assign w[973] = 16'b1000011110110001; 
assign w[974] = 16'b0001011000100110; 
assign w[975] = 16'b1100010101011000; 
assign w[976] = 16'b1011101100011001; 
assign w[977] = 16'b0110001101101100; 
assign w[978] = 16'b0111010110001111; 
assign w[979] = 16'b1011001000010110; 
assign w[980] = 16'b0100011011001001; 
assign w[981] = 16'b0101100100111011; 
assign w[982] = 16'b0010100101100101; 
assign w[983] = 16'b0110110010110101; 
assign w[984] = 16'b1001011110110011; 
assign w[985] = 16'b0001011001100110; 
assign w[986] = 16'b1100110101011001; 
assign w[987] = 16'b1011101100111001; 
assign w[988] = 16'b0110011101101100; 
assign w[989] = 16'b1111010110011111; 
assign w[990] = 16'b1011010000010110; 
assign w[991] = 16'b1000011011010001; 
assign w[992] = 16'b0101101000111011; 
assign w[993] = 16'b0100100101101001; 
assign w[994] = 16'b0110110100110101; 
assign w[995] = 16'b1010011110110101; 
assign w[996] = 16'b0001011010100110; 
assign w[997] = 16'b1101010101011010; 
assign w[998] = 16'b1011101101011001; 
assign w[999] = 16'b0110101101101101; 
assign w[1000] = 16'b0111010110101111; 
assign w[1001] = 16'b1011011000010110; 
assign w[1002] = 16'b1100011011011001; 
assign w[1003] = 16'b0101101100111011; 
assign w[1004] = 16'b0110100101101101; 
assign w[1005] = 16'b0110110110110101; 
assign w[1006] = 16'b1011011110110111; 
assign w[1007] = 16'b0001011011100110; 
assign w[1008] = 16'b1101110101011011; 
assign w[1009] = 16'b1011101101111001; 
assign w[1010] = 16'b0110111101101101; 
assign w[1011] = 16'b1111010110111111; 
assign w[1012] = 16'b1011100000010111; 
assign w[1013] = 16'b0000011011100001; 
assign w[1014] = 16'b0101110000111011; 
assign w[1015] = 16'b1000100101110001; 
assign w[1016] = 16'b0110111000110101; 
assign w[1017] = 16'b1100011110111001; 
assign w[1018] = 16'b0001011100100110; 
assign w[1019] = 16'b1110010101011100; 
assign w[1020] = 16'b1011101110011001; 
assign w[1021] = 16'b0111001101101110; 
assign w[1022] = 16'b0111010111001111; 
assign w[1023] = 16'b1011101000010111; 
assign w[1024] = 16'b0100011011101001; 
assign w[1025] = 16'b0101110100111011; 
assign w[1026] = 16'b1010100101110101; 
assign w[1027] = 16'b0110111010110101; 
assign w[1028] = 16'b1101011110111011; 
assign w[1029] = 16'b0001011101100110; 
assign w[1030] = 16'b1110110101011101; 
assign w[1031] = 16'b1011101110111001; 
assign w[1032] = 16'b0111011101101110; 
assign w[1033] = 16'b1111010111011111; 
assign w[1034] = 16'b1011110000010111; 
assign w[1035] = 16'b1000011011110001; 
assign w[1036] = 16'b0101111000111011; 
assign w[1037] = 16'b1100100101111001; 
assign w[1038] = 16'b0110111100110101; 
assign w[1039] = 16'b1110011110111101; 
assign w[1040] = 16'b0001011110100110; 
assign w[1041] = 16'b1111010101011110; 
assign w[1042] = 16'b1011101111011001; 
assign w[1043] = 16'b0111101101101111; 
assign w[1044] = 16'b0111010111101111; 
assign w[1045] = 16'b1011111000010111; 
assign w[1046] = 16'b1100011011111001; 
assign w[1047] = 16'b0101111100111011; 
assign w[1048] = 16'b1110100101111101; 
assign w[1049] = 16'b0110111110110101; 
assign w[1050] = 16'b1111011110111111; 
assign w[1051] = 16'b0001011111100110; 
assign w[1052] = 16'b1111110101011111; 
assign w[1053] = 16'b1011101111111001; 
assign w[1054] = 16'b0111111101101111; 
assign w[1055] = 16'b1111010111111111; 
assign w[1056] = 16'b1100000000011000; 
assign w[1057] = 16'b0000011100000001; 
assign w[1058] = 16'b0110000000111100; 
assign w[1059] = 16'b0000100110000001; 
assign w[1060] = 16'b0111000000110110; 
assign w[1061] = 16'b0000011111000001; 
assign w[1062] = 16'b0001100000100111; 
assign w[1063] = 16'b0000010101100000; 
assign w[1064] = 16'b1011110000011001; 
assign w[1065] = 16'b1000001101110000; 
assign w[1066] = 16'b0111011000001111; 
assign w[1067] = 16'b1100001000011000; 
assign w[1068] = 16'b0100011100001001; 
assign w[1069] = 16'b0110000100111100; 
assign w[1070] = 16'b0010100110000101; 
assign w[1071] = 16'b0111000010110110; 
assign w[1072] = 16'b0001011111000011; 
assign w[1073] = 16'b0001100001100111; 
assign w[1074] = 16'b0000110101100001; 
assign w[1075] = 16'b1011110000111001; 
assign w[1076] = 16'b1000011101110000; 
assign w[1077] = 16'b1111011000011111; 
assign w[1078] = 16'b1100010000011000; 
assign w[1079] = 16'b1000011100010001; 
assign w[1080] = 16'b0110001000111100; 
assign w[1081] = 16'b0100100110001001; 
assign w[1082] = 16'b0111000100110110; 
assign w[1083] = 16'b0010011111000101; 
assign w[1084] = 16'b0001100010100111; 
assign w[1085] = 16'b0001010101100010; 
assign w[1086] = 16'b1011110001011001; 
assign w[1087] = 16'b1000101101110001; 
assign w[1088] = 16'b0111011000101111; 
assign w[1089] = 16'b1100011000011000; 
assign w[1090] = 16'b1100011100011001; 
assign w[1091] = 16'b0110001100111100; 
assign w[1092] = 16'b0110100110001101; 
assign w[1093] = 16'b0111000110110110; 
assign w[1094] = 16'b0011011111000111; 
assign w[1095] = 16'b0001100011100111; 
assign w[1096] = 16'b0001110101100011; 
assign w[1097] = 16'b1011110001111001; 
assign w[1098] = 16'b1000111101110001; 
assign w[1099] = 16'b1111011000111111; 
assign w[1100] = 16'b1100100000011001; 
assign w[1101] = 16'b0000011100100001; 
assign w[1102] = 16'b0110010000111100; 
assign w[1103] = 16'b1000100110010001; 
assign w[1104] = 16'b0111001000110110; 
assign w[1105] = 16'b0100011111001001; 
assign w[1106] = 16'b0001100100100111; 
assign w[1107] = 16'b0010010101100100; 
assign w[1108] = 16'b1011110010011001; 
assign w[1109] = 16'b1001001101110010; 
assign w[1110] = 16'b0111011001001111; 
assign w[1111] = 16'b1100101000011001; 
assign w[1112] = 16'b0100011100101001; 
assign w[1113] = 16'b0110010100111100; 
assign w[1114] = 16'b1010100110010101; 
assign w[1115] = 16'b0111001010110110; 
assign w[1116] = 16'b0101011111001011; 
assign w[1117] = 16'b0001100101100111; 
assign w[1118] = 16'b0010110101100101; 
assign w[1119] = 16'b1011110010111001; 
assign w[1120] = 16'b1001011101110010; 
assign w[1121] = 16'b1111011001011111; 
assign w[1122] = 16'b1100110000011001; 
assign w[1123] = 16'b1000011100110001; 
assign w[1124] = 16'b0110011000111100; 
assign w[1125] = 16'b1100100110011001; 
assign w[1126] = 16'b0111001100110110; 
assign w[1127] = 16'b0110011111001101; 
assign w[1128] = 16'b0001100110100111; 
assign w[1129] = 16'b0011010101100110; 
assign w[1130] = 16'b1011110011011001; 
assign w[1131] = 16'b1001101101110011; 
assign w[1132] = 16'b0111011001101111; 
assign w[1133] = 16'b1100111000011001; 
assign w[1134] = 16'b1100011100111001; 
assign w[1135] = 16'b0110011100111100; 
assign w[1136] = 16'b1110100110011101; 
assign w[1137] = 16'b0111001110110110; 
assign w[1138] = 16'b0111011111001111; 
assign w[1139] = 16'b0001100111100111; 
assign w[1140] = 16'b0011110101100111; 
assign w[1141] = 16'b1011110011111001; 
assign w[1142] = 16'b1001111101110011; 
assign w[1143] = 16'b1111011001111111; 
assign w[1144] = 16'b1101000000011010; 
assign w[1145] = 16'b0000011101000001; 
assign w[1146] = 16'b0110100000111101; 
assign w[1147] = 16'b0000100110100001; 
assign w[1148] = 16'b0111010000110110; 
assign w[1149] = 16'b1000011111010001; 
assign w[1150] = 16'b0001101000100111; 
assign w[1151] = 16'b0100010101101000; 
assign w[1152] = 16'b1011110100011001; 
assign w[1153] = 16'b1010001101110100; 
assign w[1154] = 16'b0111011010001111; 
assign w[1155] = 16'b1101001000011010; 
assign w[1156] = 16'b0100011101001001; 
assign w[1157] = 16'b0110100100111101; 
assign w[1158] = 16'b0010100110100101; 
assign w[1159] = 16'b0111010010110110; 
assign w[1160] = 16'b1001011111010011; 
assign w[1161] = 16'b0001101001100111; 
assign w[1162] = 16'b0100110101101001; 
assign w[1163] = 16'b1011110100111001; 
assign w[1164] = 16'b1010011101110100; 
assign w[1165] = 16'b1111011010011111; 
assign w[1166] = 16'b1101010000011010; 
assign w[1167] = 16'b1000011101010001; 
assign w[1168] = 16'b0110101000111101; 
assign w[1169] = 16'b0100100110101001; 
assign w[1170] = 16'b0111010100110110; 
assign w[1171] = 16'b1010011111010101; 
assign w[1172] = 16'b0001101010100111; 
assign w[1173] = 16'b0101010101101010; 
assign w[1174] = 16'b1011110101011001; 
assign w[1175] = 16'b1010101101110101; 
assign w[1176] = 16'b0111011010101111; 
assign w[1177] = 16'b1101011000011010; 
assign w[1178] = 16'b1100011101011001; 
assign w[1179] = 16'b0110101100111101; 
assign w[1180] = 16'b0110100110101101; 
assign w[1181] = 16'b0111010110110110; 
assign w[1182] = 16'b1011011111010111; 
assign w[1183] = 16'b0001101011100111; 
assign w[1184] = 16'b0101110101101011; 
assign w[1185] = 16'b1011110101111001; 
assign w[1186] = 16'b1010111101110101; 
assign w[1187] = 16'b1111011010111111; 
assign w[1188] = 16'b1101100000011011; 
assign w[1189] = 16'b0000011101100001; 
assign w[1190] = 16'b0110110000111101; 
assign w[1191] = 16'b1000100110110001; 
assign w[1192] = 16'b0111011000110110; 
assign w[1193] = 16'b1100011111011001; 
assign w[1194] = 16'b0001101100100111; 
assign w[1195] = 16'b0110010101101100; 
assign w[1196] = 16'b1011110110011001; 
assign w[1197] = 16'b1011001101110110; 
assign w[1198] = 16'b0111011011001111; 
assign w[1199] = 16'b1101101000011011; 
assign w[1200] = 16'b0100011101101001; 
assign w[1201] = 16'b0110110100111101; 
assign w[1202] = 16'b1010100110110101; 
assign w[1203] = 16'b0111011010110110; 
assign w[1204] = 16'b1101011111011011; 
assign w[1205] = 16'b0001101101100111; 
assign w[1206] = 16'b0110110101101101; 
assign w[1207] = 16'b1011110110111001; 
assign w[1208] = 16'b1011011101110110; 
assign w[1209] = 16'b1111011011011111; 
assign w[1210] = 16'b1101110000011011; 
assign w[1211] = 16'b1000011101110001; 
assign w[1212] = 16'b0110111000111101; 
assign w[1213] = 16'b1100100110111001; 
assign w[1214] = 16'b0111011100110110; 
assign w[1215] = 16'b1110011111011101; 
assign w[1216] = 16'b0001101110100111; 
assign w[1217] = 16'b0111010101101110; 
assign w[1218] = 16'b1011110111011001; 
assign w[1219] = 16'b1011101101110111; 
assign w[1220] = 16'b0111011011101111; 
assign w[1221] = 16'b1101111000011011; 
assign w[1222] = 16'b1100011101111001; 
assign w[1223] = 16'b0110111100111101; 
assign w[1224] = 16'b1110100110111101; 
assign w[1225] = 16'b0111011110110110; 
assign w[1226] = 16'b1111011111011111; 
assign w[1227] = 16'b0001101111100111; 
assign w[1228] = 16'b0111110101101111; 
assign w[1229] = 16'b1011110111111001; 
assign w[1230] = 16'b1011111101110111; 
assign w[1231] = 16'b1111011011111111; 
assign w[1232] = 16'b1110000000011100; 
assign w[1233] = 16'b0000011110000001; 
assign w[1234] = 16'b0111000000111110; 
assign w[1235] = 16'b0000100111000001; 
assign w[1236] = 16'b0111100000110111; 
assign w[1237] = 16'b0000011111100001; 
assign w[1238] = 16'b0001110000100111; 
assign w[1239] = 16'b1000010101110000; 
assign w[1240] = 16'b1011111000011001; 
assign w[1241] = 16'b1100001101111000; 
assign w[1242] = 16'b0111011100001111; 
assign w[1243] = 16'b1110001000011100; 
assign w[1244] = 16'b0100011110001001; 
assign w[1245] = 16'b0111000100111110; 
assign w[1246] = 16'b0010100111000101; 
assign w[1247] = 16'b0111100010110111; 
assign w[1248] = 16'b0001011111100011; 
assign w[1249] = 16'b0001110001100111; 
assign w[1250] = 16'b1000110101110001; 
assign w[1251] = 16'b1011111000111001; 
assign w[1252] = 16'b1100011101111000; 
assign w[1253] = 16'b1111011100011111; 
assign w[1254] = 16'b1110010000011100; 
assign w[1255] = 16'b1000011110010001; 
assign w[1256] = 16'b0111001000111110; 
assign w[1257] = 16'b0100100111001001; 
assign w[1258] = 16'b0111100100110111; 
assign w[1259] = 16'b0010011111100101; 
assign w[1260] = 16'b0001110010100111; 
assign w[1261] = 16'b1001010101110010; 
assign w[1262] = 16'b1011111001011001; 
assign w[1263] = 16'b1100101101111001; 
assign w[1264] = 16'b0111011100101111; 
assign w[1265] = 16'b1110011000011100; 
assign w[1266] = 16'b1100011110011001; 
assign w[1267] = 16'b0111001100111110; 
assign w[1268] = 16'b0110100111001101; 
assign w[1269] = 16'b0111100110110111; 
assign w[1270] = 16'b0011011111100111; 
assign w[1271] = 16'b0001110011100111; 
assign w[1272] = 16'b1001110101110011; 
assign w[1273] = 16'b1011111001111001; 
assign w[1274] = 16'b1100111101111001; 
assign w[1275] = 16'b1111011100111111; 
assign w[1276] = 16'b1110100000011101; 
assign w[1277] = 16'b0000011110100001; 
assign w[1278] = 16'b0111010000111110; 
assign w[1279] = 16'b1000100111010001; 
assign w[1280] = 16'b0111101000110111; 
assign w[1281] = 16'b0100011111101001; 
assign w[1282] = 16'b0001110100100111; 
assign w[1283] = 16'b1010010101110100; 
assign w[1284] = 16'b1011111010011001; 
assign w[1285] = 16'b1101001101111010; 
assign w[1286] = 16'b0111011101001111; 
assign w[1287] = 16'b1110101000011101; 
assign w[1288] = 16'b0100011110101001; 
assign w[1289] = 16'b0111010100111110; 
assign w[1290] = 16'b1010100111010101; 
assign w[1291] = 16'b0111101010110111; 
assign w[1292] = 16'b0101011111101011; 
assign w[1293] = 16'b0001110101100111; 
assign w[1294] = 16'b1010110101110101; 
assign w[1295] = 16'b1011111010111001; 
assign w[1296] = 16'b1101011101111010; 
assign w[1297] = 16'b1111011101011111; 
assign w[1298] = 16'b1110110000011101; 
assign w[1299] = 16'b1000011110110001; 
assign w[1300] = 16'b0111011000111110; 
assign w[1301] = 16'b1100100111011001; 
assign w[1302] = 16'b0111101100110111; 
assign w[1303] = 16'b0110011111101101; 
assign w[1304] = 16'b0001110110100111; 
assign w[1305] = 16'b1011010101110110; 
assign w[1306] = 16'b1011111011011001; 
assign w[1307] = 16'b1101101101111011; 
assign w[1308] = 16'b0111011101101111; 
assign w[1309] = 16'b1110111000011101; 
assign w[1310] = 16'b1100011110111001; 
assign w[1311] = 16'b0111011100111110; 
assign w[1312] = 16'b1110100111011101; 
assign w[1313] = 16'b0111101110110111; 
assign w[1314] = 16'b0111011111101111; 
assign w[1315] = 16'b0001110111100111; 
assign w[1316] = 16'b1011110101110111; 
assign w[1317] = 16'b1011111011111001; 
assign w[1318] = 16'b1101111101111011; 
assign w[1319] = 16'b1111011101111111; 
assign w[1320] = 16'b1111000000011110; 
assign w[1321] = 16'b0000011111000001; 
assign w[1322] = 16'b0111100000111111; 
assign w[1323] = 16'b0000100111100001; 
assign w[1324] = 16'b0111110000110111; 
assign w[1325] = 16'b1000011111110001; 
assign w[1326] = 16'b0001111000100111; 
assign w[1327] = 16'b1100010101111000; 
assign w[1328] = 16'b1011111100011001; 
assign w[1329] = 16'b1110001101111100; 
assign w[1330] = 16'b0111011110001111; 
assign w[1331] = 16'b1111001000011110; 
assign w[1332] = 16'b0100011111001001; 
assign w[1333] = 16'b0111100100111111; 
assign w[1334] = 16'b0010100111100101; 
assign w[1335] = 16'b0111110010110111; 
assign w[1336] = 16'b1001011111110011; 
assign w[1337] = 16'b0001111001100111; 
assign w[1338] = 16'b1100110101111001; 
assign w[1339] = 16'b1011111100111001; 
assign w[1340] = 16'b1110011101111100; 
assign w[1341] = 16'b1111011110011111; 
assign w[1342] = 16'b1111010000011110; 
assign w[1343] = 16'b1000011111010001; 
assign w[1344] = 16'b0111101000111111; 
assign w[1345] = 16'b0100100111101001; 
assign w[1346] = 16'b0111110100110111; 
assign w[1347] = 16'b1010011111110101; 
assign w[1348] = 16'b0001111010100111; 
assign w[1349] = 16'b1101010101111010; 
assign w[1350] = 16'b1011111101011001; 
assign w[1351] = 16'b1110101101111101; 
assign w[1352] = 16'b0111011110101111; 
assign w[1353] = 16'b1111011000011110; 
assign w[1354] = 16'b1100011111011001; 
assign w[1355] = 16'b0111101100111111; 
assign w[1356] = 16'b0110100111101101; 
assign w[1357] = 16'b0111110110110111; 
assign w[1358] = 16'b1011011111110111; 
assign w[1359] = 16'b0001111011100111; 
assign w[1360] = 16'b1101110101111011; 
assign w[1361] = 16'b1011111101111001; 
assign w[1362] = 16'b1110111101111101; 
assign w[1363] = 16'b1111011110111111; 
assign w[1364] = 16'b1111100000011111; 
assign w[1365] = 16'b0000011111100001; 
assign w[1366] = 16'b0111110000111111; 
assign w[1367] = 16'b1000100111110001; 
assign w[1368] = 16'b0111111000110111; 
assign w[1369] = 16'b1100011111111001; 
assign w[1370] = 16'b0001111100100111; 
assign w[1371] = 16'b1110010101111100; 
assign w[1372] = 16'b1011111110011001; 
assign w[1373] = 16'b1111001101111110; 
assign w[1374] = 16'b0111011111001111; 
assign w[1375] = 16'b1111101000011111; 
assign w[1376] = 16'b0100011111101001; 
assign w[1377] = 16'b0111110100111111; 
assign w[1378] = 16'b1010100111110101; 
assign w[1379] = 16'b0111111010110111; 
assign w[1380] = 16'b1101011111111011; 
assign w[1381] = 16'b0001111101100111; 
assign w[1382] = 16'b1110110101111101; 
assign w[1383] = 16'b1011111110111001; 
assign w[1384] = 16'b1111011101111110; 
assign w[1385] = 16'b1111011111011111; 
assign w[1386] = 16'b1111110000011111; 
assign w[1387] = 16'b1000011111110001; 
assign w[1388] = 16'b0111111000111111; 
assign w[1389] = 16'b1100100111111001; 
assign w[1390] = 16'b0111111100110111; 
assign w[1391] = 16'b1110011111111101; 
assign w[1392] = 16'b0001111110100111; 
assign w[1393] = 16'b1111010101111110; 
assign w[1394] = 16'b1011111111011001; 
assign w[1395] = 16'b1111101101111111; 
assign w[1396] = 16'b0111011111101111; 
assign w[1397] = 16'b1111111000011111; 
assign w[1398] = 16'b1100011111111001; 
assign w[1399] = 16'b0111111100111111; 
assign w[1400] = 16'b1110100111111101; 
assign w[1401] = 16'b0111111110110111; 
assign w[1402] = 16'b1111011111111111; 
assign w[1403] = 16'b0001111111100111; 
assign w[1404] = 16'b1111110101111111; 
assign w[1405] = 16'b1011111111111001; 
assign w[1406] = 16'b1111111101111111; 
assign w[1407] = 16'b1111011111111110; 

initial begin
	repeat(10)@(posedge dCLK);
	repeat(100)begin
		repeat(10240) begin
			dFM = 0;
			dDAT = w[wrdCnt2][bitCnt];
			bitCnt <= bitCnt - 1'b1;
			if(bitCnt == 4'd15) begin
				wrdCnt <= wrdCnt + 1'b1;
				wrdCnt2 <= wrdCnt2 + 1'b1;
				if(wrdCnt == 5'd9) begin
					strNum <= strNum + 1'b1;
				end else
				if(wrdCnt == 5'd19) begin
					strNum <= strNum + 1'b1;
					if (strNum == 6'd63) begin
						frmNum <= frmNum + 1'b1;
						dFM = 1;
					end
					wrdCnt <= 5'b0;
				end
				if (wrdCnt2 == 10'd1407) begin
					wrdCnt2 <= 10'd0;
				end

			end
			@(posedge dCLK);
		end
	end
	$stop;
end


DTFM DTFM_tb(
	.clk(clk),
	.clk80(clk80),
	.dCLK(dCLK),
	.dFM(dFM),
	.dDAT(dDAT),
	.FRM(out)
);

endmodule

module PowerController(
	input 					clk,
	input 					reset,
	input 		[11:0] 	curr_pwr,		//0-4095
	output 		[6:0]		duty
);

endmodule

module distributor(
);

endmodule

module DTFM (
	input clk,
	input dCLK,
	input dFM,
	input dDAT,
	output FRM
);


endmodule
